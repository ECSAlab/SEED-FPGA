------------------------------------------------------------------------------------------------
--  This source is dedicated to the research paper enttled                                    --
--  "An 8-bit Serialized Architecture of SEED Block Cipher for Constrained Devices"           --
--  on IET Circuits, Devices & Systems journal                                                --
--  Authors : Lampros Pyrgas, Filippos Pirpilidis and Paris Kitsos                            --
--  Institute: University of the Peloponnese                                                  --
--  Department: Electrical and Computer Engineering                                           --
--                                                                                            --
--  This source is distributed in the hope that it will be useful, but WITHOUT ANY WARRANTY.  --
------------------------------------------------------------------------------------------------

module GF2(
input [1:0] a,
input [1:0] b,
output [1:0] ab
);

assign ab[1] = (a[1]&b[0])^(a[0]&b[1])^(a[1]&b[1]);
assign ab[0] = (a[1]&b[1])^(a[0]&b[0]);
endmodule
